module andGate(
    input D,
    input E,
    output out
    );

assign out= D & E;
endmodule