`timescale 1ns/1ns
`include "registerMemory.v"

module register_memory_tb;

initial begin

	$dumpfile("register_memory_tb.vcd");
	$dumpvars;
    
	


end
endmodule